module main

fn main() {
	if ab {
		eprintln('test')
	} else if c {
		eprintln('abc')
	} else {
		eprintln(123)
	}
}