module ast

pub struct File {
pub:
	stmts []Stmt
}