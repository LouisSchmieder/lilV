module main

import test as abc

// test
/* test */

pub fn main() {}
