module token

struct Position {
	file string
	line_nr int
	char_nr int
}