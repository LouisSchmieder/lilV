module test

fn test(test i8) int {}

['test': 123; abc]
fn main() {}
