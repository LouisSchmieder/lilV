module token

struct Position {
	file string
pub:
	line_nr int
	char_nr int
}