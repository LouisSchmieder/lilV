module main

// test
/* test */

fn main() {}
