module token

struct Position {
pub:
	file string
	line_nr int
	char_nr int
}