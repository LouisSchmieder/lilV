module main

pub const abc = 'def'

const (
	test = 123
	abc = 544
)